package trans;
 typedef struct {
    int burst_id;
    logic [7:0] data;
    logic valid;
} transaction_t;
endpackage
